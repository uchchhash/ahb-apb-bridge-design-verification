package ahb_env_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"
    
    import apb_agent_pkg::*;
    import ahb_agent_pkg::*;
    
    
    `include "def_tb.sv"
    `include "ahb_scoreboard.sv"
    `include "ahb_env_config.sv"
    `include "ahb_env.sv"

endpackage


