package ahb_seq_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"
    
    import ahb_agent_pkg::ahb_seq_item;
    
    `include "def_tb.sv"
    `include "ahb_base_sequence.sv"
    `include "ahb_reset_sequence.sv"
    `include "ahb_write_sequence.sv"
    `include "ahb_read_sequence.sv"

endpackage