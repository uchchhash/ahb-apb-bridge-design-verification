package ahb_agent_pkg;

    import uvm_pkg::*;
    `include "uvm_macros.svh"

    `include "ahb_seq_item.sv"
    
    `include "def_tb.sv"
    `include "ahb_seqr.sv"
    `include "ahb_agent_config.sv"
    `include "ahb_drv.sv"
    `include "ahb_mntr.sv"
    `include "ahb_agent.sv"

endpackage

